module TESTCASE ();
     
endmodule
