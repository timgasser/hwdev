// Include the mips1 top defines
`include "mips1_top_defines.v"

// PSX Top level defines