module TESTCASE ();


endmodule // testcase
